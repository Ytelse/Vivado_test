library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package alu_ops is

  type alu_op_t is (ALU_OP_ADD, ALU_OP_SUB, ALU_OP_LT, ALU_OP_SHIFT);

end package alu_ops;
